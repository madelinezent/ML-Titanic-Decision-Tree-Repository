// Titanic Tree
digraph {
	<__main__.DTNode object at 0x7f957ac61390> [label=Sex]
	<__main__.DTNode object at 0x7f957ac39e10> [label=Pclass]
	<__main__.DTNode object at 0x7f957ac61390> -> <__main__.DTNode object at 0x7f957ac39e10> [label=female]
	<__main__.DTNode object at 0x7f957aca9ad0> [label=Parch]
	<__main__.DTNode object at 0x7f957ac39e10> -> <__main__.DTNode object at 0x7f957aca9ad0> [label=1]
	<__main__.DTNode object at 0x7f957aca9b50> [label=alive]
	<__main__.DTNode object at 0x7f957aca9ad0> -> <__main__.DTNode object at 0x7f957aca9b50> [label=0]
	<__main__.DTNode object at 0x7f957acbc310> [label=Age]
	<__main__.DTNode object at 0x7f957aca9ad0> -> <__main__.DTNode object at 0x7f957acbc310> [label=2]
	<__main__.DTNode object at 0x7f957acbc250> [label=SibSp]
	<__main__.DTNode object at 0x7f957acbc310> -> <__main__.DTNode object at 0x7f957acbc250> [label="young adult"]
	<__main__.DTNode object at 0x7f9576c8f290> [label=alive]
	<__main__.DTNode object at 0x7f957acbc250> -> <__main__.DTNode object at 0x7f9576c8f290> [label=2]
	<__main__.DTNode object at 0x7f9576c8f190> [label=dead]
	<__main__.DTNode object at 0x7f957acbc250> -> <__main__.DTNode object at 0x7f9576c8f190> [label=1]
	<__main__.DTNode object at 0x7f957aca9810> [label=alive]
	<__main__.DTNode object at 0x7f957acbc310> -> <__main__.DTNode object at 0x7f957aca9810> [label="middle-aged"]
	<__main__.DTNode object at 0x7f957acbc810> [label=alive]
	<__main__.DTNode object at 0x7f957acbc310> -> <__main__.DTNode object at 0x7f957acbc810> [label=teen]
	<__main__.DTNode object at 0x7f957ac9fd10> [label=alive]
	<__main__.DTNode object at 0x7f957aca9ad0> -> <__main__.DTNode object at 0x7f957ac9fd10> [label=1]
	<__main__.DTNode object at 0x7f957aca9b10> [label=Age]
	<__main__.DTNode object at 0x7f957ac39e10> -> <__main__.DTNode object at 0x7f957aca9b10> [label=2]
	<__main__.DTNode object at 0x7f957acbc0d0> [label=alive]
	<__main__.DTNode object at 0x7f957aca9b10> -> <__main__.DTNode object at 0x7f957acbc0d0> [label=teen]
	<__main__.DTNode object at 0x7f9576c8fa10> [label=alive]
	<__main__.DTNode object at 0x7f957aca9b10> -> <__main__.DTNode object at 0x7f9576c8fa10> [label=child]
	<__main__.DTNode object at 0x7f957aca9b90> [label=SibSp]
	<__main__.DTNode object at 0x7f957aca9b10> -> <__main__.DTNode object at 0x7f957aca9b90> [label="young adult"]
	<__main__.DTNode object at 0x7f957acbc550> [label=alive]
	<__main__.DTNode object at 0x7f957aca9b90> -> <__main__.DTNode object at 0x7f957acbc550> [label=2]
	<__main__.DTNode object at 0x7f957acbc490> [label=alive]
	<__main__.DTNode object at 0x7f957aca9b90> -> <__main__.DTNode object at 0x7f957acbc490> [label=0]
	<__main__.DTNode object at 0x7f957afbc9d0> [label=alive]
	<__main__.DTNode object at 0x7f957aca9b90> -> <__main__.DTNode object at 0x7f957afbc9d0> [label=3]
	<__main__.DTNode object at 0x7f957ad12910> [label=Embarked]
	<__main__.DTNode object at 0x7f957aca9b90> -> <__main__.DTNode object at 0x7f957ad12910> [label=1]
	<__main__.DTNode object at 0x7f95788100d0> [label=dead]
	<__main__.DTNode object at 0x7f957ad12910> -> <__main__.DTNode object at 0x7f95788100d0> [label=S]
	<__main__.DTNode object at 0x7f957ad12190> [label=alive]
	<__main__.DTNode object at 0x7f957ad12910> -> <__main__.DTNode object at 0x7f957ad12190> [label=C]
	<__main__.DTNode object at 0x7f9576c8f0d0> [label=alive]
	<__main__.DTNode object at 0x7f957aca9b10> -> <__main__.DTNode object at 0x7f9576c8f0d0> [label="middle-aged"]
	<__main__.DTNode object at 0x7f957aca9ed0> [label=dead]
	<__main__.DTNode object at 0x7f957aca9b10> -> <__main__.DTNode object at 0x7f957aca9ed0> [label=old]
	<__main__.DTNode object at 0x7f957aca9f90> [label=Fare]
	<__main__.DTNode object at 0x7f957ac39e10> -> <__main__.DTNode object at 0x7f957aca9f90> [label=3]
	<__main__.DTNode object at 0x7f957afbce90> [label=Age]
	<__main__.DTNode object at 0x7f957aca9f90> -> <__main__.DTNode object at 0x7f957afbce90> [label="lower class"]
	<__main__.DTNode object at 0x7f957ad127d0> [label=Parch]
	<__main__.DTNode object at 0x7f957afbce90> -> <__main__.DTNode object at 0x7f957ad127d0> [label="young adult"]
	<__main__.DTNode object at 0x7f957ad12410> [label=dead]
	<__main__.DTNode object at 0x7f957ad127d0> -> <__main__.DTNode object at 0x7f957ad12410> [label=0]
	<__main__.DTNode object at 0x7f957ad12dd0> [label=alive]
	<__main__.DTNode object at 0x7f957ad127d0> -> <__main__.DTNode object at 0x7f957ad12dd0> [label=2]
	<__main__.DTNode object at 0x7f957ad125d0> [label=dead]
	<__main__.DTNode object at 0x7f957afbce90> -> <__main__.DTNode object at 0x7f957ad125d0> [label=child]
	<__main__.DTNode object at 0x7f957ad12d10> [label=alive]
	<__main__.DTNode object at 0x7f957afbce90> -> <__main__.DTNode object at 0x7f957ad12d10> [label="middle-aged"]
	<__main__.DTNode object at 0x7f957acbc650> [label=SibSp]
	<__main__.DTNode object at 0x7f957aca9f90> -> <__main__.DTNode object at 0x7f957acbc650> [label="middle class"]
	<__main__.DTNode object at 0x7f957afbc710> [label=Parch]
	<__main__.DTNode object at 0x7f957acbc650> -> <__main__.DTNode object at 0x7f957afbc710> [label=1]
	<__main__.DTNode object at 0x7f957ad12c10> [label=dead]
	<__main__.DTNode object at 0x7f957afbc710> -> <__main__.DTNode object at 0x7f957ad12c10> [label=0]
	<__main__.DTNode object at 0x7f957ad12d90> [label=dead]
	<__main__.DTNode object at 0x7f957afbc710> -> <__main__.DTNode object at 0x7f957ad12d90> [label=1]
	<__main__.DTNode object at 0x7f957ad12810> [label=dead]
	<__main__.DTNode object at 0x7f957afbc710> -> <__main__.DTNode object at 0x7f957ad12810> [label=2]
	<__main__.DTNode object at 0x7f957ad12e10> [label=Age]
	<__main__.DTNode object at 0x7f957acbc650> -> <__main__.DTNode object at 0x7f957ad12e10> [label=0]
	<__main__.DTNode object at 0x7f957ad126d0> [label=alive]
	<__main__.DTNode object at 0x7f957ad12e10> -> <__main__.DTNode object at 0x7f957ad126d0> [label="young adult"]
	<__main__.DTNode object at 0x7f957ad12a50> [label=dead]
	<__main__.DTNode object at 0x7f957ad12e10> -> <__main__.DTNode object at 0x7f957ad12a50> [label=teen]
	<__main__.DTNode object at 0x7f957ad12e90> [label=dead]
	<__main__.DTNode object at 0x7f957ad12e10> -> <__main__.DTNode object at 0x7f957ad12e90> [label="middle-aged"]
	<__main__.DTNode object at 0x7f957ad12b10> [label=alive]
	<__main__.DTNode object at 0x7f957ad12e10> -> <__main__.DTNode object at 0x7f957ad12b10> [label=child]
	<__main__.DTNode object at 0x7f957acbc2d0> [label=alive]
	<__main__.DTNode object at 0x7f957acbc650> -> <__main__.DTNode object at 0x7f957acbc2d0> [label=2]
	<__main__.DTNode object at 0x7f957ad122d0> [label=Age]
	<__main__.DTNode object at 0x7f957acbc650> -> <__main__.DTNode object at 0x7f957ad122d0> [label=3]
	<__main__.DTNode object at 0x7f957ad12ed0> [label=alive]
	<__main__.DTNode object at 0x7f957ad122d0> -> <__main__.DTNode object at 0x7f957ad12ed0> [label="middle-aged"]
	<__main__.DTNode object at 0x7f957ad12710> [label=dead]
	<__main__.DTNode object at 0x7f957ad122d0> -> <__main__.DTNode object at 0x7f957ad12710> [label=child]
	<__main__.DTNode object at 0x7f957acbc510> [label=SibSp]
	<__main__.DTNode object at 0x7f957aca9f90> -> <__main__.DTNode object at 0x7f957acbc510> [label=poor]
	<__main__.DTNode object at 0x7f957ad12f90> [label=Parch]
	<__main__.DTNode object at 0x7f957acbc510> -> <__main__.DTNode object at 0x7f957ad12f90> [label=0]
	<__main__.DTNode object at 0x7f957ad12b90> [label=alive]
	<__main__.DTNode object at 0x7f957ad12f90> -> <__main__.DTNode object at 0x7f957ad12b90> [label=0]
	<__main__.DTNode object at 0x7f957ad12150> [label=dead]
	<__main__.DTNode object at 0x7f957ad12f90> -> <__main__.DTNode object at 0x7f957ad12150> [label=2]
	<__main__.DTNode object at 0x7f957ad12f10> [label=dead]
	<__main__.DTNode object at 0x7f957acbc510> -> <__main__.DTNode object at 0x7f957ad12f10> [label=1]
	<__main__.DTNode object at 0x7f957ad12bd0> [label=Age]
	<__main__.DTNode object at 0x7f957aca9f90> -> <__main__.DTNode object at 0x7f957ad12bd0> [label="upper class"]
	<__main__.DTNode object at 0x7f957ad12990> [label=dead]
	<__main__.DTNode object at 0x7f957ad12bd0> -> <__main__.DTNode object at 0x7f957ad12990> [label="middle-aged"]
	<__main__.DTNode object at 0x7f957ad12cd0> [label=SibSp]
	<__main__.DTNode object at 0x7f957ad12bd0> -> <__main__.DTNode object at 0x7f957ad12cd0> [label=child]
	<__main__.DTNode object at 0x7f957ad096d0> [label=dead]
	<__main__.DTNode object at 0x7f957ad12cd0> -> <__main__.DTNode object at 0x7f957ad096d0> [label=4]
	<__main__.DTNode object at 0x7f957ad12ad0> [label=dead]
	<__main__.DTNode object at 0x7f957ad12bd0> -> <__main__.DTNode object at 0x7f957ad12ad0> [label="young adult"]
	<__main__.DTNode object at 0x7f9576cb60d0> [label=Fare]
	<__main__.DTNode object at 0x7f957ac61390> -> <__main__.DTNode object at 0x7f9576cb60d0> [label=male]
	<__main__.DTNode object at 0x7f957afbc310> [label=Embarked]
	<__main__.DTNode object at 0x7f9576cb60d0> -> <__main__.DTNode object at 0x7f957afbc310> [label=poor]
	<__main__.DTNode object at 0x7f957acbcdd0> [label=Age]
	<__main__.DTNode object at 0x7f957afbc310> -> <__main__.DTNode object at 0x7f957acbcdd0> [label=S]
	<__main__.DTNode object at 0x7f957ad09350> [label=SibSp]
	<__main__.DTNode object at 0x7f957acbcdd0> -> <__main__.DTNode object at 0x7f957ad09350> [label="young adult"]
	<__main__.DTNode object at 0x7f957ad09b50> [label=dead]
	<__main__.DTNode object at 0x7f957ad09350> -> <__main__.DTNode object at 0x7f957ad09b50> [label=0]
	<__main__.DTNode object at 0x7f957ad09250> [label=dead]
	<__main__.DTNode object at 0x7f957ad09350> -> <__main__.DTNode object at 0x7f957ad09250> [label=1]
	<__main__.DTNode object at 0x7f957ad12a90> [label=Pclass]
	<__main__.DTNode object at 0x7f957acbcdd0> -> <__main__.DTNode object at 0x7f957ad12a90> [label="middle-aged"]
	<__main__.DTNode object at 0x7f957ad09290> [label=dead]
	<__main__.DTNode object at 0x7f957ad12a90> -> <__main__.DTNode object at 0x7f957ad09290> [label=3]
	<__main__.DTNode object at 0x7f957ad09650> [label=dead]
	<__main__.DTNode object at 0x7f957ad12a90> -> <__main__.DTNode object at 0x7f957ad09650> [label=1]
	<__main__.DTNode object at 0x7f957ad124d0> [label=dead]
	<__main__.DTNode object at 0x7f957acbcdd0> -> <__main__.DTNode object at 0x7f957ad124d0> [label=old]
	<__main__.DTNode object at 0x7f957ad12950> [label=dead]
	<__main__.DTNode object at 0x7f957acbcdd0> -> <__main__.DTNode object at 0x7f957ad12950> [label=teen]
	<__main__.DTNode object at 0x7f957ad12550> [label=Age]
	<__main__.DTNode object at 0x7f957afbc310> -> <__main__.DTNode object at 0x7f957ad12550> [label=Q]
	<__main__.DTNode object at 0x7f957ad12850> [label=dead]
	<__main__.DTNode object at 0x7f957ad12550> -> <__main__.DTNode object at 0x7f957ad12850> [label="middle-aged"]
	<__main__.DTNode object at 0x7f957ad12f50> [label=Pclass]
	<__main__.DTNode object at 0x7f957ad12550> -> <__main__.DTNode object at 0x7f957ad12f50> [label="young adult"]
	<__main__.DTNode object at 0x7f957ad09850> [label=dead]
	<__main__.DTNode object at 0x7f957ad12f50> -> <__main__.DTNode object at 0x7f957ad09850> [label=3]
	<__main__.DTNode object at 0x7f957acbc690> [label=dead]
	<__main__.DTNode object at 0x7f957afbc310> -> <__main__.DTNode object at 0x7f957acbc690> [label=C]
	<__main__.DTNode object at 0x7f957ac39ed0> [label=Pclass]
	<__main__.DTNode object at 0x7f9576cb60d0> -> <__main__.DTNode object at 0x7f957ac39ed0> [label="middle class"]
	<__main__.DTNode object at 0x7f957ad123d0> [label=Age]
	<__main__.DTNode object at 0x7f957ac39ed0> -> <__main__.DTNode object at 0x7f957ad123d0> [label=2]
	<__main__.DTNode object at 0x7f957ad09d50> [label=SibSp]
	<__main__.DTNode object at 0x7f957ad123d0> -> <__main__.DTNode object at 0x7f957ad09d50> [label="middle-aged"]
	<__main__.DTNode object at 0x7f957ad09610> [label=dead]
	<__main__.DTNode object at 0x7f957ad09d50> -> <__main__.DTNode object at 0x7f957ad09610> [label=0]
	<__main__.DTNode object at 0x7f957ad09b90> [label=dead]
	<__main__.DTNode object at 0x7f957ad09d50> -> <__main__.DTNode object at 0x7f957ad09b90> [label=1]
	<__main__.DTNode object at 0x7f957afbc290> [label=Embarked]
	<__main__.DTNode object at 0x7f957ad123d0> -> <__main__.DTNode object at 0x7f957afbc290> [label="young adult"]
	<__main__.DTNode object at 0x7f957ad09e50> [label=dead]
	<__main__.DTNode object at 0x7f957afbc290> -> <__main__.DTNode object at 0x7f957ad09e50> [label=S]
	<__main__.DTNode object at 0x7f957ad09590> [label=dead]
	<__main__.DTNode object at 0x7f957afbc290> -> <__main__.DTNode object at 0x7f957ad09590> [label=C]
	<__main__.DTNode object at 0x7f957ad09f50> [label=dead]
	<__main__.DTNode object at 0x7f957ad123d0> -> <__main__.DTNode object at 0x7f957ad09f50> [label=teen]
	<__main__.DTNode object at 0x7f957ad097d0> [label=alive]
	<__main__.DTNode object at 0x7f957ad123d0> -> <__main__.DTNode object at 0x7f957ad097d0> [label=child]
	<__main__.DTNode object at 0x7f957acbc050> [label=Age]
	<__main__.DTNode object at 0x7f957ac39ed0> -> <__main__.DTNode object at 0x7f957acbc050> [label=1]
	<__main__.DTNode object at 0x7f957ad09710> [label=Embarked]
	<__main__.DTNode object at 0x7f957acbc050> -> <__main__.DTNode object at 0x7f957ad09710> [label="young adult"]
	<__main__.DTNode object at 0x7f957ad09110> [label=alive]
	<__main__.DTNode object at 0x7f957ad09710> -> <__main__.DTNode object at 0x7f957ad09110> [label=S]
	<__main__.DTNode object at 0x7f957ad09cd0> [label=dead]
	<__main__.DTNode object at 0x7f957ad09710> -> <__main__.DTNode object at 0x7f957ad09cd0> [label=C]
	<__main__.DTNode object at 0x7f957ad12790> [label=SibSp]
	<__main__.DTNode object at 0x7f957acbc050> -> <__main__.DTNode object at 0x7f957ad12790> [label="middle-aged"]
	<__main__.DTNode object at 0x7f957ad093d0> [label=dead]
	<__main__.DTNode object at 0x7f957ad12790> -> <__main__.DTNode object at 0x7f957ad093d0> [label=0]
	<__main__.DTNode object at 0x7f957ad12b50> [label=dead]
	<__main__.DTNode object at 0x7f957acbc050> -> <__main__.DTNode object at 0x7f957ad12b50> [label=old]
	<__main__.DTNode object at 0x7f957afbc110> [label=Embarked]
	<__main__.DTNode object at 0x7f957ac39ed0> -> <__main__.DTNode object at 0x7f957afbc110> [label=3]
	<__main__.DTNode object at 0x7f957ad09c50> [label=dead]
	<__main__.DTNode object at 0x7f957afbc110> -> <__main__.DTNode object at 0x7f957ad09c50> [label=S]
	<__main__.DTNode object at 0x7f957aca97d0> [label=Parch]
	<__main__.DTNode object at 0x7f957afbc110> -> <__main__.DTNode object at 0x7f957aca97d0> [label=C]
	<__main__.DTNode object at 0x7f957ad09c90> [label=dead]
	<__main__.DTNode object at 0x7f957aca97d0> -> <__main__.DTNode object at 0x7f957ad09c90> [label=0]
	<__main__.DTNode object at 0x7f957ad09c10> [label=alive]
	<__main__.DTNode object at 0x7f957aca97d0> -> <__main__.DTNode object at 0x7f957ad09c10> [label=1]
	<__main__.DTNode object at 0x7f957ad09510> [label=SibSp]
	<__main__.DTNode object at 0x7f957afbc110> -> <__main__.DTNode object at 0x7f957ad09510> [label=Q]
	<__main__.DTNode object at 0x7f957ad09fd0> [label=dead]
	<__main__.DTNode object at 0x7f957ad09510> -> <__main__.DTNode object at 0x7f957ad09fd0> [label=4]
	<__main__.DTNode object at 0x7f957ad09790> [label=alive]
	<__main__.DTNode object at 0x7f957ad09510> -> <__main__.DTNode object at 0x7f957ad09790> [label=2]
	<__main__.DTNode object at 0x7f957ad09690> [label=dead]
	<__main__.DTNode object at 0x7f957ad09510> -> <__main__.DTNode object at 0x7f957ad09690> [label=1]
	<__main__.DTNode object at 0x7f957acbc7d0> [label=Age]
	<__main__.DTNode object at 0x7f9576cb60d0> -> <__main__.DTNode object at 0x7f957acbc7d0> [label=rich]
	<__main__.DTNode object at 0x7f957ad09e90> [label=Pclass]
	<__main__.DTNode object at 0x7f957acbc7d0> -> <__main__.DTNode object at 0x7f957ad09e90> [label="young adult"]
	<__main__.DTNode object at 0x7f957ad09750> [label=SibSp]
	<__main__.DTNode object at 0x7f957ad09e90> -> <__main__.DTNode object at 0x7f957ad09750> [label=1]
	<__main__.DTNode object at 0x7f957ad095d0> [label=dead]
	<__main__.DTNode object at 0x7f957ad09750> -> <__main__.DTNode object at 0x7f957ad095d0> [label=1]
	<__main__.DTNode object at 0x7f957afbc4d0> [label=SibSp]
	<__main__.DTNode object at 0x7f957acbc7d0> -> <__main__.DTNode object at 0x7f957afbc4d0> [label="middle-aged"]
	<__main__.DTNode object at 0x7f957ad09f10> [label=alive]
	<__main__.DTNode object at 0x7f957afbc4d0> -> <__main__.DTNode object at 0x7f957ad09f10> [label=0]
	<__main__.DTNode object at 0x7f957ad09050> [label=alive]
	<__main__.DTNode object at 0x7f957afbc4d0> -> <__main__.DTNode object at 0x7f957ad09050> [label=1]
	<__main__.DTNode object at 0x7f957ad09dd0> [label=dead]
	<__main__.DTNode object at 0x7f957afbc4d0> -> <__main__.DTNode object at 0x7f957ad09dd0> [label=2]
	<__main__.DTNode object at 0x7f957ad12650> [label=dead]
	<__main__.DTNode object at 0x7f957acbc7d0> -> <__main__.DTNode object at 0x7f957ad12650> [label=old]
	<__main__.DTNode object at 0x7f957a4b08d0> [label=alive]
	<__main__.DTNode object at 0x7f957acbc7d0> -> <__main__.DTNode object at 0x7f957a4b08d0> [label=teen]
	<__main__.DTNode object at 0x7f957ad091d0> [label=alive]
	<__main__.DTNode object at 0x7f957acbc7d0> -> <__main__.DTNode object at 0x7f957ad091d0> [label=child]
	<__main__.DTNode object at 0x7f957ad12690> [label=SibSp]
	<__main__.DTNode object at 0x7f9576cb60d0> -> <__main__.DTNode object at 0x7f957ad12690> [label="upper class"]
	<__main__.DTNode object at 0x7f957ad09bd0> [label=Pclass]
	<__main__.DTNode object at 0x7f957ad12690> -> <__main__.DTNode object at 0x7f957ad09bd0> [label=0]
	<__main__.DTNode object at 0x7f957ad09950> [label=Age]
	<__main__.DTNode object at 0x7f957ad09bd0> -> <__main__.DTNode object at 0x7f957ad09950> [label=1]
	<__main__.DTNode object at 0x7f957ad09a50> [label=dead]
	<__main__.DTNode object at 0x7f957ad09950> -> <__main__.DTNode object at 0x7f957ad09a50> [label=old]
	<__main__.DTNode object at 0x7f957ad297d0> [label=alive]
	<__main__.DTNode object at 0x7f957ad09950> -> <__main__.DTNode object at 0x7f957ad297d0> [label="young adult"]
	<__main__.DTNode object at 0x7f957ad29510> [label=dead]
	<__main__.DTNode object at 0x7f957ad09950> -> <__main__.DTNode object at 0x7f957ad29510> [label="middle-aged"]
	<__main__.DTNode object at 0x7f957ad29150> [label=dead]
	<__main__.DTNode object at 0x7f957ad09950> -> <__main__.DTNode object at 0x7f957ad29150> [label=elderly]
	<__main__.DTNode object at 0x7f957ad090d0> [label=Age]
	<__main__.DTNode object at 0x7f957ad09bd0> -> <__main__.DTNode object at 0x7f957ad090d0> [label=2]
	<__main__.DTNode object at 0x7f957ad29890> [label=dead]
	<__main__.DTNode object at 0x7f957ad090d0> -> <__main__.DTNode object at 0x7f957ad29890> [label=teen]
	<__main__.DTNode object at 0x7f957ad09d90> [label=alive]
	<__main__.DTNode object at 0x7f957ad090d0> -> <__main__.DTNode object at 0x7f957ad09d90> [label=child]
	<__main__.DTNode object at 0x7f957ad29610> [label=dead]
	<__main__.DTNode object at 0x7f957ad090d0> -> <__main__.DTNode object at 0x7f957ad29610> [label="young adult"]
	<__main__.DTNode object at 0x7f957ad09910> [label=alive]
	<__main__.DTNode object at 0x7f957ad09bd0> -> <__main__.DTNode object at 0x7f957ad09910> [label=3]
	<__main__.DTNode object at 0x7f957ad09150> [label=Age]
	<__main__.DTNode object at 0x7f957ad12690> -> <__main__.DTNode object at 0x7f957ad09150> [label=1]
	<__main__.DTNode object at 0x7f957ad09890> [label=Embarked]
	<__main__.DTNode object at 0x7f957ad09150> -> <__main__.DTNode object at 0x7f957ad09890> [label="young adult"]
	<__main__.DTNode object at 0x7f957ad29d10> [label=alive]
	<__main__.DTNode object at 0x7f957ad09890> -> <__main__.DTNode object at 0x7f957ad29d10> [label=C]
	<__main__.DTNode object at 0x7f957ad299d0> [label=dead]
	<__main__.DTNode object at 0x7f957ad09890> -> <__main__.DTNode object at 0x7f957ad299d0> [label=S]
	<__main__.DTNode object at 0x7f957ad098d0> [label=Pclass]
	<__main__.DTNode object at 0x7f957ad09150> -> <__main__.DTNode object at 0x7f957ad098d0> [label="middle-aged"]
	<__main__.DTNode object at 0x7f957ad29e50> [label=dead]
	<__main__.DTNode object at 0x7f957ad098d0> -> <__main__.DTNode object at 0x7f957ad29e50> [label=3]
	<__main__.DTNode object at 0x7f957ad12e50> [label=dead]
	<__main__.DTNode object at 0x7f957ad098d0> -> <__main__.DTNode object at 0x7f957ad12e50> [label=2]
	<__main__.DTNode object at 0x7f957ad29710> [label=dead]
	<__main__.DTNode object at 0x7f957ad098d0> -> <__main__.DTNode object at 0x7f957ad29710> [label=1]
	<__main__.DTNode object at 0x7f957ad09190> [label=dead]
	<__main__.DTNode object at 0x7f957ad09150> -> <__main__.DTNode object at 0x7f957ad09190> [label=old]
	<__main__.DTNode object at 0x7f957acbc4d0> [label=dead]
	<__main__.DTNode object at 0x7f957ad12690> -> <__main__.DTNode object at 0x7f957acbc4d0> [label=5]
	<__main__.DTNode object at 0x7f957ad092d0> [label=dead]
	<__main__.DTNode object at 0x7f957ad12690> -> <__main__.DTNode object at 0x7f957ad092d0> [label=4]
	<__main__.DTNode object at 0x7f957ad09390> [label=dead]
	<__main__.DTNode object at 0x7f957ad12690> -> <__main__.DTNode object at 0x7f957ad09390> [label=8]
	<__main__.DTNode object at 0x7f957ad09450> [label=dead]
	<__main__.DTNode object at 0x7f957ad12690> -> <__main__.DTNode object at 0x7f957ad09450> [label=2]
	<__main__.DTNode object at 0x7f957acca750> [label=Age]
	<__main__.DTNode object at 0x7f9576cb60d0> -> <__main__.DTNode object at 0x7f957acca750> [label="lower class"]
	<__main__.DTNode object at 0x7f957ad09490> [label=Pclass]
	<__main__.DTNode object at 0x7f957acca750> -> <__main__.DTNode object at 0x7f957ad09490> [label="young adult"]
	<__main__.DTNode object at 0x7f957ad291d0> [label=SibSp]
	<__main__.DTNode object at 0x7f957ad09490> -> <__main__.DTNode object at 0x7f957ad291d0> [label=3]
	<__main__.DTNode object at 0x7f957ad29790> [label=dead]
	<__main__.DTNode object at 0x7f957ad291d0> -> <__main__.DTNode object at 0x7f957ad29790> [label=0]
	<__main__.DTNode object at 0x7f957ad29b10> [label=dead]
	<__main__.DTNode object at 0x7f957ad291d0> -> <__main__.DTNode object at 0x7f957ad29b10> [label=2]
	<__main__.DTNode object at 0x7f957ad29490> [label=dead]
	<__main__.DTNode object at 0x7f957ad09490> -> <__main__.DTNode object at 0x7f957ad29490> [label=2]
	<__main__.DTNode object at 0x7f957ad09090> [label=dead]
	<__main__.DTNode object at 0x7f957acca750> -> <__main__.DTNode object at 0x7f957ad09090> [label=teen]
	<__main__.DTNode object at 0x7f957ad09d10> [label=dead]
	<__main__.DTNode object at 0x7f957acca750> -> <__main__.DTNode object at 0x7f957ad09d10> [label="middle-aged"]
	<__main__.DTNode object at 0x7f957ad09550> [label=alive]
	<__main__.DTNode object at 0x7f957acca750> -> <__main__.DTNode object at 0x7f957ad09550> [label=old]
	<__main__.DTNode object at 0x7f957ad09e10> [label=alive]
	<__main__.DTNode object at 0x7f957acca750> -> <__main__.DTNode object at 0x7f957ad09e10> [label=child]
}
