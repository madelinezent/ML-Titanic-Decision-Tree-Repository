// Titanic Tree
digraph {
	<__main__.DTNode object at 0x7f8254743790> [label=Sex]
	<__main__.DTNode object at 0x7f82513d6410> [label=Pclass]
	<__main__.DTNode object at 0x7f8254743790> -> <__main__.DTNode object at 0x7f82513d6410> [label=female]
	<__main__.DTNode object at 0x7f8253bd1650> [label=Parch]
	<__main__.DTNode object at 0x7f82513d6410> -> <__main__.DTNode object at 0x7f8253bd1650> [label=1]
	<__main__.DTNode object at 0x7f825494ec50> [label=alive]
	<__main__.DTNode object at 0x7f8253bd1650> -> <__main__.DTNode object at 0x7f825494ec50> [label=0]
	<__main__.DTNode object at 0x7f82548f5a50> [label=Age]
	<__main__.DTNode object at 0x7f8253bd1650> -> <__main__.DTNode object at 0x7f82548f5a50> [label=2]
	<__main__.DTNode object at 0x7f82549182d0> [label=SibSp]
	<__main__.DTNode object at 0x7f82548f5a50> -> <__main__.DTNode object at 0x7f82549182d0> [label="young adult"]
	<__main__.DTNode object at 0x7f8254918350> [label=alive]
	<__main__.DTNode object at 0x7f82549182d0> -> <__main__.DTNode object at 0x7f8254918350> [label=2]
	<__main__.DTNode object at 0x7f8254918150> [label=dead]
	<__main__.DTNode object at 0x7f82549182d0> -> <__main__.DTNode object at 0x7f8254918150> [label=1]
	<__main__.DTNode object at 0x7f82514fa190> [label=alive]
	<__main__.DTNode object at 0x7f82548f5a50> -> <__main__.DTNode object at 0x7f82514fa190> [label="middle-aged"]
	<__main__.DTNode object at 0x7f82514fa390> [label=alive]
	<__main__.DTNode object at 0x7f82548f5a50> -> <__main__.DTNode object at 0x7f82514fa390> [label=teen]
	<__main__.DTNode object at 0x7f82514fa490> [label=alive]
	<__main__.DTNode object at 0x7f8253bd1650> -> <__main__.DTNode object at 0x7f82514fa490> [label=1]
	<__main__.DTNode object at 0x7f825473c150> [label=Age]
	<__main__.DTNode object at 0x7f82513d6410> -> <__main__.DTNode object at 0x7f825473c150> [label=2]
	<__main__.DTNode object at 0x7f82548fdad0> [label=alive]
	<__main__.DTNode object at 0x7f825473c150> -> <__main__.DTNode object at 0x7f82548fdad0> [label=teen]
	<__main__.DTNode object at 0x7f824f355710> [label=alive]
	<__main__.DTNode object at 0x7f825473c150> -> <__main__.DTNode object at 0x7f824f355710> [label=child]
	<__main__.DTNode object at 0x7f825494e210> [label=SibSp]
	<__main__.DTNode object at 0x7f825473c150> -> <__main__.DTNode object at 0x7f825494e210> [label="young adult"]
	<__main__.DTNode object at 0x7f82548fded0> [label=alive]
	<__main__.DTNode object at 0x7f825494e210> -> <__main__.DTNode object at 0x7f82548fded0> [label=2]
	<__main__.DTNode object at 0x7f82548fdf90> [label=alive]
	<__main__.DTNode object at 0x7f825494e210> -> <__main__.DTNode object at 0x7f82548fdf90> [label=0]
	<__main__.DTNode object at 0x7f82548fda10> [label=alive]
	<__main__.DTNode object at 0x7f825494e210> -> <__main__.DTNode object at 0x7f82548fda10> [label=3]
	<__main__.DTNode object at 0x7f8254bf9f90> [label=Embarked]
	<__main__.DTNode object at 0x7f825494e210> -> <__main__.DTNode object at 0x7f8254bf9f90> [label=1]
	<__main__.DTNode object at 0x7f8254bf9950> [label=dead]
	<__main__.DTNode object at 0x7f8254bf9f90> -> <__main__.DTNode object at 0x7f8254bf9950> [label=S]
	<__main__.DTNode object at 0x7f8254bf9c90> [label=alive]
	<__main__.DTNode object at 0x7f8254bf9f90> -> <__main__.DTNode object at 0x7f8254bf9c90> [label=C]
	<__main__.DTNode object at 0x7f82549092d0> [label=alive]
	<__main__.DTNode object at 0x7f825473c150> -> <__main__.DTNode object at 0x7f82549092d0> [label="middle-aged"]
	<__main__.DTNode object at 0x7f82548edd90> [label=dead]
	<__main__.DTNode object at 0x7f825473c150> -> <__main__.DTNode object at 0x7f82548edd90> [label=old]
	<__main__.DTNode object at 0x7f8254918390> [label=Fare]
	<__main__.DTNode object at 0x7f82513d6410> -> <__main__.DTNode object at 0x7f8254918390> [label=3]
	<__main__.DTNode object at 0x7f82548fdd50> [label=Age]
	<__main__.DTNode object at 0x7f8254918390> -> <__main__.DTNode object at 0x7f82548fdd50> [label="lower class"]
	<__main__.DTNode object at 0x7f825494e150> [label=Parch]
	<__main__.DTNode object at 0x7f82548fdd50> -> <__main__.DTNode object at 0x7f825494e150> [label="young adult"]
	<__main__.DTNode object at 0x7f82549489d0> [label=dead]
	<__main__.DTNode object at 0x7f825494e150> -> <__main__.DTNode object at 0x7f82549489d0> [label=0]
	<__main__.DTNode object at 0x7f825494e590> [label=alive]
	<__main__.DTNode object at 0x7f825494e150> -> <__main__.DTNode object at 0x7f825494e590> [label=2]
	<__main__.DTNode object at 0x7f8254bf9cd0> [label=dead]
	<__main__.DTNode object at 0x7f82548fdd50> -> <__main__.DTNode object at 0x7f8254bf9cd0> [label=child]
	<__main__.DTNode object at 0x7f825494ea50> [label=alive]
	<__main__.DTNode object at 0x7f82548fdd50> -> <__main__.DTNode object at 0x7f825494ea50> [label="middle-aged"]
	<__main__.DTNode object at 0x7f8254bf9e90> [label=SibSp]
	<__main__.DTNode object at 0x7f8254918390> -> <__main__.DTNode object at 0x7f8254bf9e90> [label="middle class"]
	<__main__.DTNode object at 0x7f825494ef10> [label=Parch]
	<__main__.DTNode object at 0x7f8254bf9e90> -> <__main__.DTNode object at 0x7f825494ef10> [label=1]
	<__main__.DTNode object at 0x7f8254bf9f10> [label=dead]
	<__main__.DTNode object at 0x7f825494ef10> -> <__main__.DTNode object at 0x7f8254bf9f10> [label=0]
	<__main__.DTNode object at 0x7f8254948610> [label=dead]
	<__main__.DTNode object at 0x7f825494ef10> -> <__main__.DTNode object at 0x7f8254948610> [label=1]
	<__main__.DTNode object at 0x7f8254948090> [label=dead]
	<__main__.DTNode object at 0x7f825494ef10> -> <__main__.DTNode object at 0x7f8254948090> [label=2]
	<__main__.DTNode object at 0x7f82548fdb10> [label=Age]
	<__main__.DTNode object at 0x7f8254bf9e90> -> <__main__.DTNode object at 0x7f82548fdb10> [label=0]
	<__main__.DTNode object at 0x7f8254948e10> [label=alive]
	<__main__.DTNode object at 0x7f82548fdb10> -> <__main__.DTNode object at 0x7f8254948e10> [label="young adult"]
	<__main__.DTNode object at 0x7f825494ef50> [label=dead]
	<__main__.DTNode object at 0x7f82548fdb10> -> <__main__.DTNode object at 0x7f825494ef50> [label=teen]
	<__main__.DTNode object at 0x7f825494e290> [label=dead]
	<__main__.DTNode object at 0x7f82548fdb10> -> <__main__.DTNode object at 0x7f825494e290> [label="middle-aged"]
	<__main__.DTNode object at 0x7f82549480d0> [label=alive]
	<__main__.DTNode object at 0x7f82548fdb10> -> <__main__.DTNode object at 0x7f82549480d0> [label=child]
	<__main__.DTNode object at 0x7f8254918250> [label=alive]
	<__main__.DTNode object at 0x7f8254bf9e90> -> <__main__.DTNode object at 0x7f8254918250> [label=2]
	<__main__.DTNode object at 0x7f825494e910> [label=Age]
	<__main__.DTNode object at 0x7f8254bf9e90> -> <__main__.DTNode object at 0x7f825494e910> [label=3]
	<__main__.DTNode object at 0x7f8254948890> [label=alive]
	<__main__.DTNode object at 0x7f825494e910> -> <__main__.DTNode object at 0x7f8254948890> [label="middle-aged"]
	<__main__.DTNode object at 0x7f8254948d50> [label=dead]
	<__main__.DTNode object at 0x7f825494e910> -> <__main__.DTNode object at 0x7f8254948d50> [label=child]
	<__main__.DTNode object at 0x7f825494eed0> [label=SibSp]
	<__main__.DTNode object at 0x7f8254918390> -> <__main__.DTNode object at 0x7f825494eed0> [label=poor]
	<__main__.DTNode object at 0x7f8254bf9450> [label=Parch]
	<__main__.DTNode object at 0x7f825494eed0> -> <__main__.DTNode object at 0x7f8254bf9450> [label=0]
	<__main__.DTNode object at 0x7f8254948b50> [label=alive]
	<__main__.DTNode object at 0x7f8254bf9450> -> <__main__.DTNode object at 0x7f8254948b50> [label=0]
	<__main__.DTNode object at 0x7f82549486d0> [label=dead]
	<__main__.DTNode object at 0x7f8254bf9450> -> <__main__.DTNode object at 0x7f82549486d0> [label=2]
	<__main__.DTNode object at 0x7f8254bf99d0> [label=dead]
	<__main__.DTNode object at 0x7f825494eed0> -> <__main__.DTNode object at 0x7f8254bf99d0> [label=1]
	<__main__.DTNode object at 0x7f8254918210> [label=Age]
	<__main__.DTNode object at 0x7f8254918390> -> <__main__.DTNode object at 0x7f8254918210> [label="upper class"]
	<__main__.DTNode object at 0x7f8254948510> [label=dead]
	<__main__.DTNode object at 0x7f8254918210> -> <__main__.DTNode object at 0x7f8254948510> [label="middle-aged"]
	<__main__.DTNode object at 0x7f825494e550> [label=SibSp]
	<__main__.DTNode object at 0x7f8254918210> -> <__main__.DTNode object at 0x7f825494e550> [label=child]
	<__main__.DTNode object at 0x7f8254948a90> [label=dead]
	<__main__.DTNode object at 0x7f825494e550> -> <__main__.DTNode object at 0x7f8254948a90> [label=4]
	<__main__.DTNode object at 0x7f825494e490> [label=dead]
	<__main__.DTNode object at 0x7f8254918210> -> <__main__.DTNode object at 0x7f825494e490> [label="young adult"]
	<__main__.DTNode object at 0x7f82548f5490> [label=Fare]
	<__main__.DTNode object at 0x7f8254743790> -> <__main__.DTNode object at 0x7f82548f5490> [label=male]
	<__main__.DTNode object at 0x7f8254bf9dd0> [label=Embarked]
	<__main__.DTNode object at 0x7f82548f5490> -> <__main__.DTNode object at 0x7f8254bf9dd0> [label=poor]
	<__main__.DTNode object at 0x7f8254918310> [label=Age]
	<__main__.DTNode object at 0x7f8254bf9dd0> -> <__main__.DTNode object at 0x7f8254918310> [label=S]
	<__main__.DTNode object at 0x7f8254948d90> [label=SibSp]
	<__main__.DTNode object at 0x7f8254918310> -> <__main__.DTNode object at 0x7f8254948d90> [label="young adult"]
	<__main__.DTNode object at 0x7f8254948c90> [label=dead]
	<__main__.DTNode object at 0x7f8254948d90> -> <__main__.DTNode object at 0x7f8254948c90> [label=0]
	<__main__.DTNode object at 0x7f8254948f90> [label=dead]
	<__main__.DTNode object at 0x7f8254948d90> -> <__main__.DTNode object at 0x7f8254948f90> [label=1]
	<__main__.DTNode object at 0x7f825494e390> [label=Pclass]
	<__main__.DTNode object at 0x7f8254918310> -> <__main__.DTNode object at 0x7f825494e390> [label="middle-aged"]
	<__main__.DTNode object at 0x7f8254948e90> [label=dead]
	<__main__.DTNode object at 0x7f825494e390> -> <__main__.DTNode object at 0x7f8254948e90> [label=3]
	<__main__.DTNode object at 0x7f8254948c10> [label=dead]
	<__main__.DTNode object at 0x7f825494e390> -> <__main__.DTNode object at 0x7f8254948c10> [label=1]
	<__main__.DTNode object at 0x7f825494e250> [label=dead]
	<__main__.DTNode object at 0x7f8254918310> -> <__main__.DTNode object at 0x7f825494e250> [label=old]
	<__main__.DTNode object at 0x7f8254948d10> [label=dead]
	<__main__.DTNode object at 0x7f8254918310> -> <__main__.DTNode object at 0x7f8254948d10> [label=teen]
	<__main__.DTNode object at 0x7f825494ef90> [label=Age]
	<__main__.DTNode object at 0x7f8254bf9dd0> -> <__main__.DTNode object at 0x7f825494ef90> [label=Q]
	<__main__.DTNode object at 0x7f8254948290> [label=dead]
	<__main__.DTNode object at 0x7f825494ef90> -> <__main__.DTNode object at 0x7f8254948290> [label="middle-aged"]
	<__main__.DTNode object at 0x7f82549482d0> [label=Pclass]
	<__main__.DTNode object at 0x7f825494ef90> -> <__main__.DTNode object at 0x7f82549482d0> [label="young adult"]
	<__main__.DTNode object at 0x7f8254948810> [label=dead]
	<__main__.DTNode object at 0x7f82549482d0> -> <__main__.DTNode object at 0x7f8254948810> [label=3]
	<__main__.DTNode object at 0x7f8254bf9bd0> [label=dead]
	<__main__.DTNode object at 0x7f8254bf9dd0> -> <__main__.DTNode object at 0x7f8254bf9bd0> [label=C]
	<__main__.DTNode object at 0x7f8254bf9a50> [label=Pclass]
	<__main__.DTNode object at 0x7f82548f5490> -> <__main__.DTNode object at 0x7f8254bf9a50> [label="middle class"]
	<__main__.DTNode object at 0x7f825494ec90> [label=Age]
	<__main__.DTNode object at 0x7f8254bf9a50> -> <__main__.DTNode object at 0x7f825494ec90> [label=2]
	<__main__.DTNode object at 0x7f8254948f10> [label=SibSp]
	<__main__.DTNode object at 0x7f825494ec90> -> <__main__.DTNode object at 0x7f8254948f10> [label="middle-aged"]
	<__main__.DTNode object at 0x7f8254948550> [label=dead]
	<__main__.DTNode object at 0x7f8254948f10> -> <__main__.DTNode object at 0x7f8254948550> [label=0]
	<__main__.DTNode object at 0x7f8254948a50> [label=dead]
	<__main__.DTNode object at 0x7f8254948f10> -> <__main__.DTNode object at 0x7f8254948a50> [label=1]
	<__main__.DTNode object at 0x7f8254948250> [label=Embarked]
	<__main__.DTNode object at 0x7f825494ec90> -> <__main__.DTNode object at 0x7f8254948250> [label="young adult"]
	<__main__.DTNode object at 0x7f8254948690> [label=dead]
	<__main__.DTNode object at 0x7f8254948250> -> <__main__.DTNode object at 0x7f8254948690> [label=S]
	<__main__.DTNode object at 0x7f8254948910> [label=dead]
	<__main__.DTNode object at 0x7f8254948250> -> <__main__.DTNode object at 0x7f8254948910> [label=C]
	<__main__.DTNode object at 0x7f8254948c50> [label=dead]
	<__main__.DTNode object at 0x7f825494ec90> -> <__main__.DTNode object at 0x7f8254948c50> [label=teen]
	<__main__.DTNode object at 0x7f8254948990> [label=alive]
	<__main__.DTNode object at 0x7f825494ec90> -> <__main__.DTNode object at 0x7f8254948990> [label=child]
	<__main__.DTNode object at 0x7f82541dd9d0> [label=Age]
	<__main__.DTNode object at 0x7f8254bf9a50> -> <__main__.DTNode object at 0x7f82541dd9d0> [label=1]
	<__main__.DTNode object at 0x7f8254948cd0> [label=Embarked]
	<__main__.DTNode object at 0x7f82541dd9d0> -> <__main__.DTNode object at 0x7f8254948cd0> [label="young adult"]
	<__main__.DTNode object at 0x7f8254973090> [label=alive]
	<__main__.DTNode object at 0x7f8254948cd0> -> <__main__.DTNode object at 0x7f8254973090> [label=S]
	<__main__.DTNode object at 0x7f8254948dd0> [label=dead]
	<__main__.DTNode object at 0x7f8254948cd0> -> <__main__.DTNode object at 0x7f8254948dd0> [label=C]
	<__main__.DTNode object at 0x7f8254948950> [label=SibSp]
	<__main__.DTNode object at 0x7f82541dd9d0> -> <__main__.DTNode object at 0x7f8254948950> [label="middle-aged"]
	<__main__.DTNode object at 0x7f8254948150> [label=dead]
	<__main__.DTNode object at 0x7f8254948950> -> <__main__.DTNode object at 0x7f8254948150> [label=0]
	<__main__.DTNode object at 0x7f8254948f50> [label=dead]
	<__main__.DTNode object at 0x7f82541dd9d0> -> <__main__.DTNode object at 0x7f8254948f50> [label=old]
	<__main__.DTNode object at 0x7f825494e3d0> [label=Embarked]
	<__main__.DTNode object at 0x7f8254bf9a50> -> <__main__.DTNode object at 0x7f825494e3d0> [label=3]
	<__main__.DTNode object at 0x7f8254948a10> [label=dead]
	<__main__.DTNode object at 0x7f825494e3d0> -> <__main__.DTNode object at 0x7f8254948a10> [label=S]
	<__main__.DTNode object at 0x7f8254948ed0> [label=Parch]
	<__main__.DTNode object at 0x7f825494e3d0> -> <__main__.DTNode object at 0x7f8254948ed0> [label=C]
	<__main__.DTNode object at 0x7f8254973810> [label=dead]
	<__main__.DTNode object at 0x7f8254948ed0> -> <__main__.DTNode object at 0x7f8254973810> [label=0]
	<__main__.DTNode object at 0x7f8254948490> [label=alive]
	<__main__.DTNode object at 0x7f8254948ed0> -> <__main__.DTNode object at 0x7f8254948490> [label=1]
	<__main__.DTNode object at 0x7f82549481d0> [label=SibSp]
	<__main__.DTNode object at 0x7f825494e3d0> -> <__main__.DTNode object at 0x7f82549481d0> [label=Q]
	<__main__.DTNode object at 0x7f8254973b90> [label=dead]
	<__main__.DTNode object at 0x7f82549481d0> -> <__main__.DTNode object at 0x7f8254973b90> [label=4]
	<__main__.DTNode object at 0x7f8254973390> [label=alive]
	<__main__.DTNode object at 0x7f82549481d0> -> <__main__.DTNode object at 0x7f8254973390> [label=2]
	<__main__.DTNode object at 0x7f8254973c50> [label=dead]
	<__main__.DTNode object at 0x7f82549481d0> -> <__main__.DTNode object at 0x7f8254973c50> [label=1]
	<__main__.DTNode object at 0x7f82549488d0> [label=Age]
	<__main__.DTNode object at 0x7f82548f5490> -> <__main__.DTNode object at 0x7f82549488d0> [label=rich]
	<__main__.DTNode object at 0x7f825494e350> [label=Pclass]
	<__main__.DTNode object at 0x7f82549488d0> -> <__main__.DTNode object at 0x7f825494e350> [label="young adult"]
	<__main__.DTNode object at 0x7f8254973910> [label=SibSp]
	<__main__.DTNode object at 0x7f825494e350> -> <__main__.DTNode object at 0x7f8254973910> [label=1]
	<__main__.DTNode object at 0x7f8254973290> [label=dead]
	<__main__.DTNode object at 0x7f8254973910> -> <__main__.DTNode object at 0x7f8254973290> [label=1]
	<__main__.DTNode object at 0x7f8254852d50> [label=SibSp]
	<__main__.DTNode object at 0x7f82549488d0> -> <__main__.DTNode object at 0x7f8254852d50> [label="middle-aged"]
	<__main__.DTNode object at 0x7f8254973550> [label=alive]
	<__main__.DTNode object at 0x7f8254852d50> -> <__main__.DTNode object at 0x7f8254973550> [label=0]
	<__main__.DTNode object at 0x7f82549487d0> [label=alive]
	<__main__.DTNode object at 0x7f8254852d50> -> <__main__.DTNode object at 0x7f82549487d0> [label=1]
	<__main__.DTNode object at 0x7f825494ee50> [label=dead]
	<__main__.DTNode object at 0x7f8254852d50> -> <__main__.DTNode object at 0x7f825494ee50> [label=2]
	<__main__.DTNode object at 0x7f8254948790> [label=dead]
	<__main__.DTNode object at 0x7f82549488d0> -> <__main__.DTNode object at 0x7f8254948790> [label=old]
	<__main__.DTNode object at 0x7f8254948850> [label=alive]
	<__main__.DTNode object at 0x7f82549488d0> -> <__main__.DTNode object at 0x7f8254948850> [label=teen]
	<__main__.DTNode object at 0x7f8254948bd0> [label=alive]
	<__main__.DTNode object at 0x7f82549488d0> -> <__main__.DTNode object at 0x7f8254948bd0> [label=child]
	<__main__.DTNode object at 0x7f8254948450> [label=SibSp]
	<__main__.DTNode object at 0x7f82548f5490> -> <__main__.DTNode object at 0x7f8254948450> [label="upper class"]
	<__main__.DTNode object at 0x7f825494e2d0> [label=Pclass]
	<__main__.DTNode object at 0x7f8254948450> -> <__main__.DTNode object at 0x7f825494e2d0> [label=0]
	<__main__.DTNode object at 0x7f8254973f90> [label=Age]
	<__main__.DTNode object at 0x7f825494e2d0> -> <__main__.DTNode object at 0x7f8254973f90> [label=1]
	<__main__.DTNode object at 0x7f8254973110> [label=dead]
	<__main__.DTNode object at 0x7f8254973f90> -> <__main__.DTNode object at 0x7f8254973110> [label=old]
	<__main__.DTNode object at 0x7f8254973b10> [label=alive]
	<__main__.DTNode object at 0x7f8254973f90> -> <__main__.DTNode object at 0x7f8254973b10> [label="young adult"]
	<__main__.DTNode object at 0x7f8254973890> [label=dead]
	<__main__.DTNode object at 0x7f8254973f90> -> <__main__.DTNode object at 0x7f8254973890> [label="middle-aged"]
	<__main__.DTNode object at 0x7f8254973bd0> [label=dead]
	<__main__.DTNode object at 0x7f8254973f90> -> <__main__.DTNode object at 0x7f8254973bd0> [label=elderly]
	<__main__.DTNode object at 0x7f8254973b50> [label=Age]
	<__main__.DTNode object at 0x7f825494e2d0> -> <__main__.DTNode object at 0x7f8254973b50> [label=2]
	<__main__.DTNode object at 0x7f82549732d0> [label=dead]
	<__main__.DTNode object at 0x7f8254973b50> -> <__main__.DTNode object at 0x7f82549732d0> [label=teen]
	<__main__.DTNode object at 0x7f8254973a50> [label=alive]
	<__main__.DTNode object at 0x7f8254973b50> -> <__main__.DTNode object at 0x7f8254973a50> [label=child]
	<__main__.DTNode object at 0x7f82549738d0> [label=dead]
	<__main__.DTNode object at 0x7f8254973b50> -> <__main__.DTNode object at 0x7f82549738d0> [label="young adult"]
	<__main__.DTNode object at 0x7f8254973690> [label=alive]
	<__main__.DTNode object at 0x7f825494e2d0> -> <__main__.DTNode object at 0x7f8254973690> [label=3]
	<__main__.DTNode object at 0x7f8254948b90> [label=Age]
	<__main__.DTNode object at 0x7f8254948450> -> <__main__.DTNode object at 0x7f8254948b90> [label=1]
	<__main__.DTNode object at 0x7f8254973790> [label=Embarked]
	<__main__.DTNode object at 0x7f8254948b90> -> <__main__.DTNode object at 0x7f8254973790> [label="young adult"]
	<__main__.DTNode object at 0x7f82549735d0> [label=alive]
	<__main__.DTNode object at 0x7f8254973790> -> <__main__.DTNode object at 0x7f82549735d0> [label=C]
	<__main__.DTNode object at 0x7f8254973c90> [label=dead]
	<__main__.DTNode object at 0x7f8254973790> -> <__main__.DTNode object at 0x7f8254973c90> [label=S]
	<__main__.DTNode object at 0x7f825494e190> [label=Pclass]
	<__main__.DTNode object at 0x7f8254948b90> -> <__main__.DTNode object at 0x7f825494e190> [label="middle-aged"]
	<__main__.DTNode object at 0x7f82549739d0> [label=dead]
	<__main__.DTNode object at 0x7f825494e190> -> <__main__.DTNode object at 0x7f82549739d0> [label=3]
	<__main__.DTNode object at 0x7f82549734d0> [label=dead]
	<__main__.DTNode object at 0x7f825494e190> -> <__main__.DTNode object at 0x7f82549734d0> [label=2]
	<__main__.DTNode object at 0x7f8254973950> [label=dead]
	<__main__.DTNode object at 0x7f825494e190> -> <__main__.DTNode object at 0x7f8254973950> [label=1]
	<__main__.DTNode object at 0x7f8254973650> [label=dead]
	<__main__.DTNode object at 0x7f8254948b90> -> <__main__.DTNode object at 0x7f8254973650> [label=old]
	<__main__.DTNode object at 0x7f82548fdb90> [label=dead]
	<__main__.DTNode object at 0x7f8254948450> -> <__main__.DTNode object at 0x7f82548fdb90> [label=5]
	<__main__.DTNode object at 0x7f8254948750> [label=dead]
	<__main__.DTNode object at 0x7f8254948450> -> <__main__.DTNode object at 0x7f8254948750> [label=4]
	<__main__.DTNode object at 0x7f8254948fd0> [label=dead]
	<__main__.DTNode object at 0x7f8254948450> -> <__main__.DTNode object at 0x7f8254948fd0> [label=8]
	<__main__.DTNode object at 0x7f8254948b10> [label=dead]
	<__main__.DTNode object at 0x7f8254948450> -> <__main__.DTNode object at 0x7f8254948b10> [label=2]
	<__main__.DTNode object at 0x7f82512e9a50> [label=Age]
	<__main__.DTNode object at 0x7f82548f5490> -> <__main__.DTNode object at 0x7f82512e9a50> [label="lower class"]
	<__main__.DTNode object at 0x7f8254973190> [label=Pclass]
	<__main__.DTNode object at 0x7f82512e9a50> -> <__main__.DTNode object at 0x7f8254973190> [label="young adult"]
	<__main__.DTNode object at 0x7f8254973510> [label=SibSp]
	<__main__.DTNode object at 0x7f8254973190> -> <__main__.DTNode object at 0x7f8254973510> [label=3]
	<__main__.DTNode object at 0x7f8254973f50> [label=dead]
	<__main__.DTNode object at 0x7f8254973510> -> <__main__.DTNode object at 0x7f8254973f50> [label=0]
	<__main__.DTNode object at 0x7f8254973490> [label=dead]
	<__main__.DTNode object at 0x7f8254973510> -> <__main__.DTNode object at 0x7f8254973490> [label=2]
	<__main__.DTNode object at 0x7f8254973990> [label=dead]
	<__main__.DTNode object at 0x7f8254973190> -> <__main__.DTNode object at 0x7f8254973990> [label=2]
	<__main__.DTNode object at 0x7f825494ecd0> [label=dead]
	<__main__.DTNode object at 0x7f82512e9a50> -> <__main__.DTNode object at 0x7f825494ecd0> [label=teen]
	<__main__.DTNode object at 0x7f825494e510> [label=dead]
	<__main__.DTNode object at 0x7f82512e9a50> -> <__main__.DTNode object at 0x7f825494e510> [label="middle-aged"]
	<__main__.DTNode object at 0x7f8254973e10> [label=alive]
	<__main__.DTNode object at 0x7f82512e9a50> -> <__main__.DTNode object at 0x7f8254973e10> [label=old]
	<__main__.DTNode object at 0x7f8254973cd0> [label=alive]
	<__main__.DTNode object at 0x7f82512e9a50> -> <__main__.DTNode object at 0x7f8254973cd0> [label=child]
}
